*** SPICE deck for cell tri_state_sim_4{lay} from library SCL-(4)
*** Created on Wed Oct 23, 2019 18:45:35
*** Last revised on Sat Oct 26, 2019 18:35:31
*** Written on Sat Oct 26, 2019 18:35:36 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT SCL-_4___tri_state_4 FROM CELL tri_state_4{lay}
.SUBCKT SCL-_4___tri_state_4 en en_ gnd in out vdd
Mnmos@9 net@219 in gnd gnd NMOS L=0.2U W=2.4U AS=3.04P AD=0.773P PS=13.4U PD=5.45U
Mnmos@10 out en net@219 gnd NMOS L=0.2U W=2.4U AS=0.773P AD=2.513P PS=5.45U PD=9.3U
Mpmos@6 net@240 in vdd vdd PMOS L=0.2U W=5.7U AS=4.735P AD=1.808P PS=19.9U PD=12.35U
Mpmos@7 out en_ net@240 vdd PMOS L=0.2U W=5.7U AS=1.808P AD=2.513P PS=12.35U PD=9.3U
.ENDS SCL-_4___tri_state_4

*** TOP LEVEL CELL: tri_state_sim_4{lay}
Xtri_stat@0 vdd gnd gnd in out vdd SCL-_4___tri_state_4

* Spice Code nodes in cell cell 'tri_state_sim_4{lay}'
vdd vdd 0 DC 3.3,
vin in 0 DC pulse 0 3.3 10n 1333.33ps 1333.33ps 10n,
cload out 0 96fF,
.tran 0 40n,
.measure tpdr 
+ TRIG v(in) VAL=1.65 FALL=1
+ TARG v(out) VAL=1.65 RISE=1
.measure tpdf 
+ TRIG v(in) VAL=1.65 RISE=1
+ TARG v(out) VAL=1.65 FALL=1
.include scmos18.txt
.END
