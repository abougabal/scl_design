*** SPICE deck for cell inverter_sim_8{lay} from library SCL-(4)
*** Created on Wed Oct 23, 2019 14:00:16
*** Last revised on Sat Oct 26, 2019 20:31:26
*** Written on Sat Oct 26, 2019 20:31:29 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT SCL-_4___inv_8 FROM CELL inv_8{lay}
.SUBCKT SCL-_4___inv_8 gnd in out vdd
Mnmos@0 out in gnd gnd NMOS L=0.2U W=2.4U AS=2.44P AD=2.288P PS=11U PD=9.25U
Mpmos@0 out in vdd vdd PMOS L=0.2U W=5.7U AS=4.085P AD=2.288P PS=17.3U PD=9.25U
.ENDS SCL-_4___inv_8

*** TOP LEVEL CELL: inverter_sim_8{lay}
Xinv_8@0 gnd in out vdd SCL-_4___inv_8

* Spice Code nodes in cell cell 'inverter_sim_8{lay}'
vdd vdd 0 DC 3.3,
vin in 0 DC pulse 0 3.3 10n 1333.33ps 1333.33ps 10n,
cload out 0 48fF,
.tran 0 40n,
.measure tpdr 
+ TRIG v(in) VAL=1.65 FALL=1
+ TARG v(out) VAL=1.65 RISE=1
.measure tpdf 
+ TRIG v(in) VAL=1.65 RISE=1
+ TARG v(out) VAL=1.65 FALL=1
.include scmos18.txt
.END
