*** SPICE deck for cell NOR1_sim{lay} from library SCL-(4)
*** Created on Sat Oct 19, 2019 15:10:35
*** Last revised on Sat Oct 26, 2019 20:23:24
*** Written on Sat Oct 26, 2019 20:23:29 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT SCL-_4___NOR3_1 FROM CELL NOR3_1{lay}
.SUBCKT SCL-_4___NOR3_1 A B C gnd NOR3 vdd
Mnmos_0 NOR3 A gnd gnd NMOS L=0.2U W=0.3U AS=0.973P AD=0.459P PS=5.017U PD=2.575U
Mnmos_1 gnd B NOR3 gnd NMOS L=0.2U W=0.3U AS=0.459P AD=0.973P PS=2.575U PD=5.017U
Mnmos_2 NOR3 C gnd gnd NMOS L=0.2U W=0.3U AS=0.973P AD=0.459P PS=5.017U PD=2.575U
Mpmos_0 vdd A net_27 vdd PMOS L=0.2U W=1.9U AS=0.57P AD=2.94P PS=2.5U PD=13.2U
Mpmos_1 net_27 B net_28 vdd PMOS L=0.2U W=1.9U AS=0.57P AD=0.57P PS=2.5U PD=2.5U
Mpmos_2 net_28 C NOR3 vdd PMOS L=0.2U W=1.9U AS=0.459P AD=0.57P PS=2.575U PD=2.5U
.ENDS SCL-_4___NOR3_1

*** TOP LEVEL CELL: NOR1_sim{lay}
XNOR3_1_2 A gnd gnd gnd NOR3 vdd SCL-_4___NOR3_1

* Spice Code nodes in cell cell 'NOR1_sim{lay}'
vdd vdd 0 DC 3.3,
vin A 0 DC pulse 0 3.3 10n 1333ps 1333ps 10n,
.tran 0 40n,
cload out 0 96fF
.measure tpd param='(tpdr+tpdf)/2'
.measure tpdr 
+ TRIG v(A) VAL=1.65 FALL=1
+ TARG v(NOR3) VAL=1.65 RISE=1
.measure tpdf 
+ TRIG v(A) VAL=1.65 RISE=1
+ TARG v(NOR3) VAL=1.65 FALL=1
.include scmos18.txt
.END
