*** SPICE deck for cell NAND3_1_lay_sim{lay} from library SCL
*** Created on Wed Oct 23, 2019 10:11:58
*** Last revised on Sat Oct 26, 2019 17:59:46
*** Written on Sat Oct 26, 2019 17:59:50 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT SCL__NAND3_1 FROM CELL NAND3_1{lay}
.SUBCKT SCL__NAND3_1 a b c gnd out vdd
Mnmos@0 net@16 a gnd gnd NMOS L=0.2U W=0.9U AS=2.83P AD=0.439P PS=13U PD=1.875U
Mnmos@1 net@1 b net@16 gnd NMOS L=0.2U W=0.9U AS=0.439P AD=0.451P PS=1.875U PD=1.95U
Mnmos@2 out c net@1 gnd NMOS L=0.2U W=0.9U AS=0.451P AD=0.471P PS=1.95U PD=2.413U
Mpmos@0 vdd a out vdd PMOS L=0.2U W=0.7U AS=0.471P AD=1.068P PS=2.413U PD=5.1U
Mpmos@1 out b vdd vdd PMOS L=0.2U W=0.7U AS=1.068P AD=0.471P PS=5.1U PD=2.413U
Mpmos@2 vdd c out vdd PMOS L=0.2U W=0.7U AS=0.471P AD=1.068P PS=2.413U PD=5.1U
.ENDS SCL__NAND3_1

*** TOP LEVEL CELL: NAND3_1_lay_sim{lay}
XNAND3_1@0 a vdd vdd gnd out vdd SCL__NAND3_1

* Spice Code nodes in cell cell 'NAND3_1_lay_sim{lay}'
vdd vdd 0 DC 3.3,
vin a 0 DC pulse 0 3.3 10n 1333.33ps 1333.33ps 10n,
cload out 0 96fF,
.tran 0 40n,
.measure tpdr 
+ TRIG v(a) VAL=1.65 FALL=1
+ TARG v(out) VAL=1.65 RISE=1
.measure tpdf 
+ TRIG v(a) VAL=1.65 RISE=1
+ TARG v(out) VAL=1.65 FALL=1
.include scmos18.txt
.END
