*** SPICE deck for cell inverter_sim{lay} from library SCL-(4)
*** Created on Fri Oct 18, 2019 21:59:56
*** Last revised on Sat Oct 26, 2019 19:54:59
*** Written on Sat Oct 26, 2019 19:55:03 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT SCL-_4___inv_1 FROM CELL inv_1{lay}
.SUBCKT SCL-_4___inv_1 gnd in out vdd
Mnmos_0 out in gnd gnd NMOS L=0.2U W=0.3U AS=1.28P AD=0.333P PS=7.2U PD=2.35U
Mpmos_0 out in vdd vdd PMOS L=0.2U W=0.7U AS=1.335P AD=0.333P PS=7.3U PD=2.35U
.ENDS SCL-_4___inv_1

*** TOP LEVEL CELL: inverter_sim{lay}
Xinv_1_0 gnd in out vdd SCL-_4___inv_1

* Spice Code nodes in cell cell 'inverter_sim{lay}'
vdd vdd 0 DC 3.3,
vin in 0 DC pulse 0 3.3 10n 0ps 0ps 10n,
.tran 0 40n,
cload out 0 96fF
.measure tpd param='(tpdr+tpdf)/2'
.measure tpdr 
+ TRIG v(in) VAL=1.65 FALL=1
+ TARG v(out) VAL=1.65 RISE=1
.measure tpdf 
+ TRIG v(in) VAL=1.65 RISE=1
+ TARG v(out) VAL=1.65 FALL=1
.include scmos18.txt
.END
