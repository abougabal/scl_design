*** SPICE deck for cell tri_state_sim_1{lay} from library SCL-(4)
*** Created on Sat Oct 26, 2019 20:51:55
*** Last revised on Sat Oct 26, 2019 21:19:12
*** Written on Sat Oct 26, 2019 21:19:16 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT SCL-_4___tri_state_1 FROM CELL tri_state_1{lay}
.SUBCKT SCL-_4___tri_state_1 en en_ gnd in out vdd
Mnmos@9 net@219 in gnd gnd NMOS L=0.2U W=0.6U AS=2.105P AD=0.225P PS=10.5U PD=1.8U
Mnmos@10 out en net@219 gnd NMOS L=0.2U W=0.6U AS=0.225P AD=0.633P PS=1.8U PD=3.3U
Mpmos@6 net@240 in vdd vdd PMOS L=0.2U W=1.4U AS=2.34P AD=0.51P PS=11U PD=3.7U
Mpmos@7 out en_ net@240 vdd PMOS L=0.2U W=1.4U AS=0.51P AD=0.633P PS=3.7U PD=3.3U
.ENDS SCL-_4___tri_state_1

*** TOP LEVEL CELL: tri_state_sim_1{lay}
Xtri_stat@0 vdd gnd gnd in out vdd SCL-_4___tri_state_1

* Spice Code nodes in cell cell 'tri_state_sim_1{lay}'
vdd vdd 0 DC 3.3,
vin in 0 DC pulse 0 3.3 10n 1333.33ps 1333.33ps 10n,
cload out 0 96fF,
.tran 0 40n,
.measure tpdr 
+ TRIG v(in) VAL=1.65 FALL=1
+ TARG v(out) VAL=1.65 RISE=1
.measure tpdf 
+ TRIG v(in) VAL=1.65 RISE=1
+ TARG v(out) VAL=1.65 FALL=1
.include scmos18.txt
.END
