*** SPICE deck for cell inverter_sim_4{lay} from library SCL-(4)
*** Created on Wed Oct 23, 2019 13:42:10
*** Last revised on Sat Oct 26, 2019 20:12:00
*** Written on Sat Oct 26, 2019 20:12:03 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT SCL-_4___inv_4 FROM CELL inv_4{lay}
.SUBCKT SCL-_4___inv_4 gnd in out vdd
Mnmos@0 out in gnd gnd NMOS L=0.2U W=1.2U AS=1.72P AD=1.103P PS=8.6U PD=5.05U
Mpmos@0 out in vdd vdd PMOS L=0.2U W=2.7U AS=2.435P AD=1.103P PS=11.3U PD=5.05U
.ENDS SCL-_4___inv_4

*** TOP LEVEL CELL: inverter_sim_4{lay}
Xinv_4@0 gnd in out vdd SCL-_4___inv_4

* Spice Code nodes in cell cell 'inverter_sim_4{lay}'
vdd vdd 0 DC 3.3,
vin in 0 DC pulse 0 3.3 10n 1333.33ps 1333.33ps 10n,
cload out 0 96fF,
.tran 0 40n,
.measure tpdr 
+ TRIG v(in) VAL=1.65 FALL=1
+ TARG v(out) VAL=1.65 RISE=1
.measure tpdf 
+ TRIG v(in) VAL=1.65 RISE=1
+ TARG v(out) VAL=1.65 FALL=1
.include scmos18.txt
.END
