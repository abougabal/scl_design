*** SPICE deck for cell inverter_sim_2{lay} from library SCL-(4)
*** Created on Wed Oct 23, 2019 13:24:46
*** Last revised on Sat Oct 26, 2019 21:20:15
*** Written on Sat Oct 26, 2019 21:20:27 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT SCL-_4___inv_2 FROM CELL inv_2{lay}
.SUBCKT SCL-_4___inv_2 gnd in out vdd
Mnmos_0 out in gnd gnd NMOS L=0.2U W=0.6U AS=1.36P AD=0.538P PS=7.4U PD=3.05U
Mpmos_0 out in vdd vdd PMOS L=0.2U W=1.3U AS=1.665P AD=0.538P PS=8.5U PD=3.05U
.ENDS SCL-_4___inv_2

*** TOP LEVEL CELL: inverter_sim_2{lay}
Xinv_2_0 gnd in out vdd SCL-_4___inv_2

* Spice Code nodes in cell cell 'inverter_sim_2{lay}'
vdd vdd 0 DC 3.3,
vin in 0 DC pulse 0 3.3 10n 667ps 667ps 10n,
.tran 0 40n,
cload out 0 96F
.measure tpd param='(tpdr+tpdf)/2'
.measure tpdr 
+ TRIG v(in) VAL=1.65 FALL=1
+ TARG v(out) VAL=1.65 RISE=1
.measure tpdf 
+ TRIG v(in) VAL=1.65 RISE=1
+ TARG v(out) VAL=1.65 FALL=1
.include scmos18.txt
.END
